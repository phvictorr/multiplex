`timescale 1ns/100ps
`include "main.v"

module main_tb;
    reg [31:0] A0, A1, A2, A3; // Entradas
    reg SEL1, SEL2; // Seletores (2, conforme o desenho)
    wire [31:0] C; // Saída

    main main1(A0, A1, A2, A3, SEL1, SEL2, C); // Instancia o módulo main
    initial begin
        $dumpfile("main_tb.vcd"); // Cria o arquivo de dump
        $dumpvars(0, main_tb); // Inicia o dump
        A0 = 32'b00000000000000000000000000000010; // 2
        A1 = 32'b00000000000000000000000000000011; // 3
        A2 = 32'b00000000000000000000000000000010; // 2
        A3 = 32'b00000000000000000000000000000011; // 3
        SEL1 = 1'b1; // 1   # Aqui é A3 = 1
        SEL2 = 1'b1; // 1
        #1
        A0 = 32'b00000000000000000000000000000010; // 2
        A1 = 32'b00000000000000000000000000000011; // 3
        A2 = 32'b00000000000000000000000000000010; // 2
        A3 = 32'b00000000000000000000000000000011; // 3
        SEL1 = 1'b1; // 1  # Aqui é A2 = 2
        SEL2 = 1'b0; // 0
        #1
        A0 = 32'b00000000000000000000000000000010; // 2
        A1 = 32'b00000000000000000000000000000011; // 3
        A2 = 32'b00000000000000000000000000000010; // 2
        A3 = 32'b00000000000000000000000000000011; // 3
        SEL1 = 1'b0; // 0  # Aqui é A1 = 1
        SEL2 = 1'b1; // 1
        #1
        A0 = 32'b00000000000000000000000000000010; // 2
        A1 = 32'b00000000000000000000000000000011; // 3
        A2 = 32'b00000000000000000000000000000010; // 2
        A3 = 32'b00000000000000000000000000000011; // 3
        SEL1 = 1'b0; // 0  # Aqui é A0 = 2
        SEL2 = 1'b0; // 0
        #1
        $finish; // para finalizar a simulação
    end
endmodule